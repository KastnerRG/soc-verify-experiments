`define R 32
`define C 64
