`define R 64
`define C 64
